** Profile: "SCHEMATIC1-DC simulation"  [ D:\SUT\Electronic 2\Pspice\elec2_project-schematic1-dc simulation.sim ] 

** Creating circuit file "elec2_project-schematic1-dc simulation.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.DC LIN V_V3 0 1m 0.00001 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\elec2_project-SCHEMATIC1.net" 


.END
